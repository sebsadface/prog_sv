module emptyBoard (
    output [15:0][15:0] GrnPixels
);

    GrnPixels[00] = 16'b1111111111111111;
    GrnPixels[01] = 16'b1000010000100001;
    GrnPixels[02] = 16'b1000010000100001;
    GrnPixels[03] = 16'b1000010000100001;
    GrnPixels[04] = 16'b1000010000100001;
    GrnPixels[05] = 16'b1111111111111111;
    GrnPixels[06] = 16'b1000010000100001;
    GrnPixels[07] = 16'b1000010000100001;
    GrnPixels[08] = 16'b1000010000100001;
    GrnPixels[09] = 16'b1000010000100001;
    GrnPixels[10] = 16'b1111111111111111;
    GrnPixels[11] = 16'b1000010000100001;
    GrnPixels[12] = 16'b1000010000100001;
    GrnPixels[13] = 16'b1000010000100001;
    GrnPixels[14] = 16'b1000010000100001;
    GrnPixels[15] = 16'b1111111111111111;

endmodule