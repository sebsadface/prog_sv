module edge_detector


endmodule // edge_detector