module user_input



endmodule // user_input